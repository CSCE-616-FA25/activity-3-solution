///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// File name   : test_lib.svh
///////////////////////////////////////////////////////////////////////////

`include "base_test.sv"
`include "mix_sequence_test.sv"
`include "agent_test.sv"